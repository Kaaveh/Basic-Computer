package States is 
	type myState is (RESET1, MEM_INIT, FINISH, FETCH1 , FETCH2, FETCH3, NOP1 , LDAC1 , LDAC2 , LDAC3, LDAC4 , LDAC5,
	STAC1, STAC2, STAC3, STAC4, STAC5, MVAC1, MOVR1, JUMP1, JUMP2, JUMP3, JMPZY1, JMPZY2, JMPZY3,
	JMPZN1, JMPZN2, JPNZY1, JPNZY2, JPNZY3, JPNZN1, JPNZN2, ADD1, SUB1, INAC1, CLAC1, AND1, OR1, XOR1, NOT1);  
end States;